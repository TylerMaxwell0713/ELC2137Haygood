module example_or(
	input a, b,
	output c
	);
	
	// c = a OR b
	or(c,a,b);	
endmodule